`timescale 1ns / 1ps
	
import lynxTypes::*;

`include "axi_macros.svh"
`include "lynx_macros.svh"

//
// Top Level - vcu118
//
module cyt_top (
 
 
	output wire        			c0_ddr4_act_n,
	output wire[16:0]  			c0_ddr4_adr,
	output wire[1:0]   			c0_ddr4_ba,
	output wire[0:0]   			c0_ddr4_bg,
	output wire[0:0]   			c0_ddr4_cke,
	output wire[0:0]   			c0_ddr4_odt,
	output wire[0:0]   			c0_ddr4_cs_n,
	output wire[0:0]   			c0_ddr4_ck_t,
	output wire[0:0]   			c0_ddr4_ck_c,
	output wire        			c0_ddr4_reset_n,
	inout  wire[7:0]   			c0_ddr4_dm_dbi_n,
	inout  wire[63:0]  			c0_ddr4_dq,
	inout  wire[7:0]   			c0_ddr4_dqs_t,
	inout  wire[7:0]   			c0_ddr4_dqs_c,
    input  wire        			c0_sys_clk_p,
	input  wire        			c0_sys_clk_n,
	output wire        			c1_ddr4_act_n,
	output wire[16:0]  			c1_ddr4_adr,
	output wire[1:0]   			c1_ddr4_ba,
	output wire[0:0]   			c1_ddr4_bg,
	output wire[0:0]   			c1_ddr4_cke,
	output wire[0:0]   			c1_ddr4_odt,
	output wire[0:0]   			c1_ddr4_cs_n,
	output wire[0:0]   			c1_ddr4_ck_t,
	output wire[0:0]   			c1_ddr4_ck_c,
	output wire        			c1_ddr4_reset_n,
	inout  wire[7:0]   			c1_ddr4_dm_dbi_n,   
	inout  wire[63:0]  			c1_ddr4_dq,
	inout  wire[7:0]   			c1_ddr4_dqs_t,
	inout  wire[7:0]   			c1_ddr4_dqs_c,
    	input  wire        		c1_sys_clk_p,
	input  wire        			c1_sys_clk_n,
	input  wire[0:0]            pcie_clk_clk_n,
	input  wire[0:0]            pcie_clk_clk_p,
	input  wire[15:0]           pcie_x16_rxn,
	input  wire[15:0]           pcie_x16_rxp,
	output wire[15:0]           pcie_x16_txn,
	output wire[15:0]           pcie_x16_txp,
	input  wire                 perst_n_nb,
	input  wire                 sys_reset_nb
);

	// Sys rst
	wire sys_reset;
	wire perst_n;
	
	// Main clk/rst
    wire uclk;
    wire [0:0] uresetn;
    wire nclk;
    wire [0:0] nresetn;
    wire pclk;
    wire [0:0] presetn;
    wire [0:0] lckresetn;
 
    wire xclk;
    wire [0:0] xresetn;
    wire aclk;
    wire [0:0] aresetn;

	// IRQ
	wire[N_REGIONS-1:0] usr_irq;

    // Static config
    AXI4L axi_cnfg_int ();
    AXI4L axi_cnfg ();

    // Application control
    AXI4L axi_ctrl_int [N_REGIONS] ();
    AXI4L axi_ctrl [N_REGIONS] ();
	
    // Application control AVX
    AXI4 #(.AXI4_DATA_BITS(AVX_DATA_BITS)) axim_ctrl_int [N_REGIONS] ();
    AXI4 #(.AXI4_DATA_BITS(AVX_DATA_BITS)) axim_ctrl [N_REGIONS] ();

    // Stream to application
    AXI4S axis_dyn_out_int [N_CHAN] ();
    AXI4S axis_dyn_out [N_CHAN] ();

    // Stream from application
    AXI4S axis_dyn_in_int [N_CHAN] ();
    AXI4S axis_dyn_in [N_CHAN] ();

    // Descriptor bypass
    dmaIntf dma_rd_req_int [N_CHAN] ();
    dmaIntf dma_rd_req [N_CHAN] ();
    dmaIntf dma_wr_req_int [N_CHAN] ();
    dmaIntf dma_wr_req [N_CHAN] ();
    xdmaIntf xdma_req_int [N_CHAN] ();
    
    // DMA Stats
    xdma_stat_t xdma_stats_0;
    xdma_stat_t xdma_stats_1;
    xdma_stat_t xdma_stats_2;
    xdma_stat_t xdma_stats_3;

    // MEM AXI mm
    AXI4 #(.AXI4_DATA_BITS(AXI_DDR_BITS)) axi_ddr_in [N_MEM_CHAN] ();
		
  // Lowspeed pins
    logic [2:0] lowspeed_ctrl_0;
    logic [2:0] lowspeed_ctrl_1;
	
	
	// ================-----------------------------------------------------------------
	// STATIC LAYER 
	// ================-----------------------------------------------------------------	
    design_static inst_int_static (
		.axi_cnfg_araddr(axi_cnfg_int.araddr),
        .axi_cnfg_arprot(axi_cnfg_int.arprot),
        .axi_cnfg_arready(axi_cnfg_int.arready),
        .axi_cnfg_arvalid(axi_cnfg_int.arvalid),
        .axi_cnfg_awaddr(axi_cnfg_int.awaddr),
        .axi_cnfg_awprot(axi_cnfg_int.awprot),
        .axi_cnfg_awready(axi_cnfg_int.awready),
        .axi_cnfg_awvalid(axi_cnfg_int.awvalid),
        .axi_cnfg_bready(axi_cnfg_int.bready),
        .axi_cnfg_bresp(axi_cnfg_int.bresp),
        .axi_cnfg_bvalid(axi_cnfg_int.bvalid),
        .axi_cnfg_rdata(axi_cnfg_int.rdata),
        .axi_cnfg_rready(axi_cnfg_int.rready),
        .axi_cnfg_rresp(axi_cnfg_int.rresp),
        .axi_cnfg_rvalid(axi_cnfg_int.rvalid),
        .axi_cnfg_wdata(axi_cnfg_int.wdata),
        .axi_cnfg_wready(axi_cnfg_int.wready),
        .axi_cnfg_wstrb(axi_cnfg_int.wstrb),
        .axi_cnfg_wvalid(axi_cnfg_int.wvalid),
        .axi_ctrl_0_araddr(axi_ctrl_int[0].araddr),
        .axi_ctrl_0_arprot(axi_ctrl_int[0].arprot),
        .axi_ctrl_0_arready(axi_ctrl_int[0].arready),
        .axi_ctrl_0_arvalid(axi_ctrl_int[0].arvalid),
        .axi_ctrl_0_awaddr(axi_ctrl_int[0].awaddr),
        .axi_ctrl_0_awprot(axi_ctrl_int[0].awprot),
        .axi_ctrl_0_awready(axi_ctrl_int[0].awready),
        .axi_ctrl_0_awvalid(axi_ctrl_int[0].awvalid),
        .axi_ctrl_0_bready(axi_ctrl_int[0].bready),
        .axi_ctrl_0_bresp(axi_ctrl_int[0].bresp),
        .axi_ctrl_0_bvalid(axi_ctrl_int[0].bvalid),
        .axi_ctrl_0_rdata(axi_ctrl_int[0].rdata),
        .axi_ctrl_0_rready(axi_ctrl_int[0].rready),
        .axi_ctrl_0_rresp(axi_ctrl_int[0].rresp),
        .axi_ctrl_0_rvalid(axi_ctrl_int[0].rvalid),
        .axi_ctrl_0_wdata(axi_ctrl_int[0].wdata),
        .axi_ctrl_0_wready(axi_ctrl_int[0].wready),
        .axi_ctrl_0_wstrb(axi_ctrl_int[0].wstrb),
        .axi_ctrl_0_wvalid(axi_ctrl_int[0].wvalid),
        .axi_ctrl_1_araddr(axi_ctrl_int[1].araddr),
        .axi_ctrl_1_arprot(axi_ctrl_int[1].arprot),
        .axi_ctrl_1_arready(axi_ctrl_int[1].arready),
        .axi_ctrl_1_arvalid(axi_ctrl_int[1].arvalid),
        .axi_ctrl_1_awaddr(axi_ctrl_int[1].awaddr),
        .axi_ctrl_1_awprot(axi_ctrl_int[1].awprot),
        .axi_ctrl_1_awready(axi_ctrl_int[1].awready),
        .axi_ctrl_1_awvalid(axi_ctrl_int[1].awvalid),
        .axi_ctrl_1_bready(axi_ctrl_int[1].bready),
        .axi_ctrl_1_bresp(axi_ctrl_int[1].bresp),
        .axi_ctrl_1_bvalid(axi_ctrl_int[1].bvalid),
        .axi_ctrl_1_rdata(axi_ctrl_int[1].rdata),
        .axi_ctrl_1_rready(axi_ctrl_int[1].rready),
        .axi_ctrl_1_rresp(axi_ctrl_int[1].rresp),
        .axi_ctrl_1_rvalid(axi_ctrl_int[1].rvalid),
        .axi_ctrl_1_wdata(axi_ctrl_int[1].wdata),
        .axi_ctrl_1_wready(axi_ctrl_int[1].wready),
        .axi_ctrl_1_wstrb(axi_ctrl_int[1].wstrb),
        .axi_ctrl_1_wvalid(axi_ctrl_int[1].wvalid),
        .axi_ctrl_2_araddr(axi_ctrl_int[2].araddr),
        .axi_ctrl_2_arprot(axi_ctrl_int[2].arprot),
        .axi_ctrl_2_arready(axi_ctrl_int[2].arready),
        .axi_ctrl_2_arvalid(axi_ctrl_int[2].arvalid),
        .axi_ctrl_2_awaddr(axi_ctrl_int[2].awaddr),
        .axi_ctrl_2_awprot(axi_ctrl_int[2].awprot),
        .axi_ctrl_2_awready(axi_ctrl_int[2].awready),
        .axi_ctrl_2_awvalid(axi_ctrl_int[2].awvalid),
        .axi_ctrl_2_bready(axi_ctrl_int[2].bready),
        .axi_ctrl_2_bresp(axi_ctrl_int[2].bresp),
        .axi_ctrl_2_bvalid(axi_ctrl_int[2].bvalid),
        .axi_ctrl_2_rdata(axi_ctrl_int[2].rdata),
        .axi_ctrl_2_rready(axi_ctrl_int[2].rready),
        .axi_ctrl_2_rresp(axi_ctrl_int[2].rresp),
        .axi_ctrl_2_rvalid(axi_ctrl_int[2].rvalid),
        .axi_ctrl_2_wdata(axi_ctrl_int[2].wdata),
        .axi_ctrl_2_wready(axi_ctrl_int[2].wready),
        .axi_ctrl_2_wstrb(axi_ctrl_int[2].wstrb),
        .axi_ctrl_2_wvalid(axi_ctrl_int[2].wvalid),
        .axi_ctrl_3_araddr(axi_ctrl_int[3].araddr),
        .axi_ctrl_3_arprot(axi_ctrl_int[3].arprot),
        .axi_ctrl_3_arready(axi_ctrl_int[3].arready),
        .axi_ctrl_3_arvalid(axi_ctrl_int[3].arvalid),
        .axi_ctrl_3_awaddr(axi_ctrl_int[3].awaddr),
        .axi_ctrl_3_awprot(axi_ctrl_int[3].awprot),
        .axi_ctrl_3_awready(axi_ctrl_int[3].awready),
        .axi_ctrl_3_awvalid(axi_ctrl_int[3].awvalid),
        .axi_ctrl_3_bready(axi_ctrl_int[3].bready),
        .axi_ctrl_3_bresp(axi_ctrl_int[3].bresp),
        .axi_ctrl_3_bvalid(axi_ctrl_int[3].bvalid),
        .axi_ctrl_3_rdata(axi_ctrl_int[3].rdata),
        .axi_ctrl_3_rready(axi_ctrl_int[3].rready),
        .axi_ctrl_3_rresp(axi_ctrl_int[3].rresp),
        .axi_ctrl_3_rvalid(axi_ctrl_int[3].rvalid),
        .axi_ctrl_3_wdata(axi_ctrl_int[3].wdata),
        .axi_ctrl_3_wready(axi_ctrl_int[3].wready),
        .axi_ctrl_3_wstrb(axi_ctrl_int[3].wstrb),
        .axi_ctrl_3_wvalid(axi_ctrl_int[3].wvalid),
        .axim_ctrl_0_araddr(axim_ctrl_int[0].araddr),
        .axim_ctrl_0_arburst(axim_ctrl_int[0].arburst),
        .axim_ctrl_0_arcache(axim_ctrl_int[0].arcache),
        .axim_ctrl_0_arlen(axim_ctrl_int[0].arlen),
        .axim_ctrl_0_arlock(axim_ctrl_int[0].arlock),
        .axim_ctrl_0_arprot(axim_ctrl_int[0].arprot),
        .axim_ctrl_0_arqos(axim_ctrl_int[0].arqos),
        .axim_ctrl_0_arready(axim_ctrl_int[0].arready),
        .axim_ctrl_0_arregion(axim_ctrl_int[0].arregion),
        .axim_ctrl_0_arsize(axim_ctrl_int[0].arsize),
        .axim_ctrl_0_arvalid(axim_ctrl_int[0].arvalid),
        .axim_ctrl_0_awaddr(axim_ctrl_int[0].awaddr),
        .axim_ctrl_0_awburst(axim_ctrl_int[0].awburst),
        .axim_ctrl_0_awcache(axim_ctrl_int[0].awcache),
        .axim_ctrl_0_awlen(axim_ctrl_int[0].awlen),
        .axim_ctrl_0_awlock(axim_ctrl_int[0].awlock),
        .axim_ctrl_0_awprot(axim_ctrl_int[0].awprot),
        .axim_ctrl_0_awqos(axim_ctrl_int[0].awqos),
        .axim_ctrl_0_awready(axim_ctrl_int[0].awready),
        .axim_ctrl_0_awregion(axim_ctrl_int[0].awregion),
        .axim_ctrl_0_awsize(axim_ctrl_int[0].awsize),
        .axim_ctrl_0_awvalid(axim_ctrl_int[0].awvalid),
        .axim_ctrl_0_bready(axim_ctrl_int[0].bready),
        .axim_ctrl_0_bresp(axim_ctrl_int[0].bresp),
        .axim_ctrl_0_bvalid(axim_ctrl_int[0].bvalid),
        .axim_ctrl_0_rdata(axim_ctrl_int[0].rdata),
        .axim_ctrl_0_rlast(axim_ctrl_int[0].rlast),
        .axim_ctrl_0_rready(axim_ctrl_int[0].rready),
        .axim_ctrl_0_rresp(axim_ctrl_int[0].rresp),
        .axim_ctrl_0_rvalid(axim_ctrl_int[0].rvalid),
        .axim_ctrl_0_wdata(axim_ctrl_int[0].wdata),
        .axim_ctrl_0_wlast(axim_ctrl_int[0].wlast),
        .axim_ctrl_0_wready(axim_ctrl_int[0].wready),
        .axim_ctrl_0_wstrb(axim_ctrl_int[0].wstrb),
        .axim_ctrl_0_wvalid(axim_ctrl_int[0].wvalid),
        .axim_ctrl_1_araddr(axim_ctrl_int[1].araddr),
        .axim_ctrl_1_arburst(axim_ctrl_int[1].arburst),
        .axim_ctrl_1_arcache(axim_ctrl_int[1].arcache),
        .axim_ctrl_1_arlen(axim_ctrl_int[1].arlen),
        .axim_ctrl_1_arlock(axim_ctrl_int[1].arlock),
        .axim_ctrl_1_arprot(axim_ctrl_int[1].arprot),
        .axim_ctrl_1_arqos(axim_ctrl_int[1].arqos),
        .axim_ctrl_1_arready(axim_ctrl_int[1].arready),
        .axim_ctrl_1_arregion(axim_ctrl_int[1].arregion),
        .axim_ctrl_1_arsize(axim_ctrl_int[1].arsize),
        .axim_ctrl_1_arvalid(axim_ctrl_int[1].arvalid),
        .axim_ctrl_1_awaddr(axim_ctrl_int[1].awaddr),
        .axim_ctrl_1_awburst(axim_ctrl_int[1].awburst),
        .axim_ctrl_1_awcache(axim_ctrl_int[1].awcache),
        .axim_ctrl_1_awlen(axim_ctrl_int[1].awlen),
        .axim_ctrl_1_awlock(axim_ctrl_int[1].awlock),
        .axim_ctrl_1_awprot(axim_ctrl_int[1].awprot),
        .axim_ctrl_1_awqos(axim_ctrl_int[1].awqos),
        .axim_ctrl_1_awready(axim_ctrl_int[1].awready),
        .axim_ctrl_1_awregion(axim_ctrl_int[1].awregion),
        .axim_ctrl_1_awsize(axim_ctrl_int[1].awsize),
        .axim_ctrl_1_awvalid(axim_ctrl_int[1].awvalid),
        .axim_ctrl_1_bready(axim_ctrl_int[1].bready),
        .axim_ctrl_1_bresp(axim_ctrl_int[1].bresp),
        .axim_ctrl_1_bvalid(axim_ctrl_int[1].bvalid),
        .axim_ctrl_1_rdata(axim_ctrl_int[1].rdata),
        .axim_ctrl_1_rlast(axim_ctrl_int[1].rlast),
        .axim_ctrl_1_rready(axim_ctrl_int[1].rready),
        .axim_ctrl_1_rresp(axim_ctrl_int[1].rresp),
        .axim_ctrl_1_rvalid(axim_ctrl_int[1].rvalid),
        .axim_ctrl_1_wdata(axim_ctrl_int[1].wdata),
        .axim_ctrl_1_wlast(axim_ctrl_int[1].wlast),
        .axim_ctrl_1_wready(axim_ctrl_int[1].wready),
        .axim_ctrl_1_wstrb(axim_ctrl_int[1].wstrb),
        .axim_ctrl_1_wvalid(axim_ctrl_int[1].wvalid),
        .axim_ctrl_2_araddr(axim_ctrl_int[2].araddr),
        .axim_ctrl_2_arburst(axim_ctrl_int[2].arburst),
        .axim_ctrl_2_arcache(axim_ctrl_int[2].arcache),
        .axim_ctrl_2_arlen(axim_ctrl_int[2].arlen),
        .axim_ctrl_2_arlock(axim_ctrl_int[2].arlock),
        .axim_ctrl_2_arprot(axim_ctrl_int[2].arprot),
        .axim_ctrl_2_arqos(axim_ctrl_int[2].arqos),
        .axim_ctrl_2_arready(axim_ctrl_int[2].arready),
        .axim_ctrl_2_arregion(axim_ctrl_int[2].arregion),
        .axim_ctrl_2_arsize(axim_ctrl_int[2].arsize),
        .axim_ctrl_2_arvalid(axim_ctrl_int[2].arvalid),
        .axim_ctrl_2_awaddr(axim_ctrl_int[2].awaddr),
        .axim_ctrl_2_awburst(axim_ctrl_int[2].awburst),
        .axim_ctrl_2_awcache(axim_ctrl_int[2].awcache),
        .axim_ctrl_2_awlen(axim_ctrl_int[2].awlen),
        .axim_ctrl_2_awlock(axim_ctrl_int[2].awlock),
        .axim_ctrl_2_awprot(axim_ctrl_int[2].awprot),
        .axim_ctrl_2_awqos(axim_ctrl_int[2].awqos),
        .axim_ctrl_2_awready(axim_ctrl_int[2].awready),
        .axim_ctrl_2_awregion(axim_ctrl_int[2].awregion),
        .axim_ctrl_2_awsize(axim_ctrl_int[2].awsize),
        .axim_ctrl_2_awvalid(axim_ctrl_int[2].awvalid),
        .axim_ctrl_2_bready(axim_ctrl_int[2].bready),
        .axim_ctrl_2_bresp(axim_ctrl_int[2].bresp),
        .axim_ctrl_2_bvalid(axim_ctrl_int[2].bvalid),
        .axim_ctrl_2_rdata(axim_ctrl_int[2].rdata),
        .axim_ctrl_2_rlast(axim_ctrl_int[2].rlast),
        .axim_ctrl_2_rready(axim_ctrl_int[2].rready),
        .axim_ctrl_2_rresp(axim_ctrl_int[2].rresp),
        .axim_ctrl_2_rvalid(axim_ctrl_int[2].rvalid),
        .axim_ctrl_2_wdata(axim_ctrl_int[2].wdata),
        .axim_ctrl_2_wlast(axim_ctrl_int[2].wlast),
        .axim_ctrl_2_wready(axim_ctrl_int[2].wready),
        .axim_ctrl_2_wstrb(axim_ctrl_int[2].wstrb),
        .axim_ctrl_2_wvalid(axim_ctrl_int[2].wvalid),
        .axim_ctrl_3_araddr(axim_ctrl_int[3].araddr),
        .axim_ctrl_3_arburst(axim_ctrl_int[3].arburst),
        .axim_ctrl_3_arcache(axim_ctrl_int[3].arcache),
        .axim_ctrl_3_arlen(axim_ctrl_int[3].arlen),
        .axim_ctrl_3_arlock(axim_ctrl_int[3].arlock),
        .axim_ctrl_3_arprot(axim_ctrl_int[3].arprot),
        .axim_ctrl_3_arqos(axim_ctrl_int[3].arqos),
        .axim_ctrl_3_arready(axim_ctrl_int[3].arready),
        .axim_ctrl_3_arregion(axim_ctrl_int[3].arregion),
        .axim_ctrl_3_arsize(axim_ctrl_int[3].arsize),
        .axim_ctrl_3_arvalid(axim_ctrl_int[3].arvalid),
        .axim_ctrl_3_awaddr(axim_ctrl_int[3].awaddr),
        .axim_ctrl_3_awburst(axim_ctrl_int[3].awburst),
        .axim_ctrl_3_awcache(axim_ctrl_int[3].awcache),
        .axim_ctrl_3_awlen(axim_ctrl_int[3].awlen),
        .axim_ctrl_3_awlock(axim_ctrl_int[3].awlock),
        .axim_ctrl_3_awprot(axim_ctrl_int[3].awprot),
        .axim_ctrl_3_awqos(axim_ctrl_int[3].awqos),
        .axim_ctrl_3_awready(axim_ctrl_int[3].awready),
        .axim_ctrl_3_awregion(axim_ctrl_int[3].awregion),
        .axim_ctrl_3_awsize(axim_ctrl_int[3].awsize),
        .axim_ctrl_3_awvalid(axim_ctrl_int[3].awvalid),
        .axim_ctrl_3_bready(axim_ctrl_int[3].bready),
        .axim_ctrl_3_bresp(axim_ctrl_int[3].bresp),
        .axim_ctrl_3_bvalid(axim_ctrl_int[3].bvalid),
        .axim_ctrl_3_rdata(axim_ctrl_int[3].rdata),
        .axim_ctrl_3_rlast(axim_ctrl_int[3].rlast),
        .axim_ctrl_3_rready(axim_ctrl_int[3].rready),
        .axim_ctrl_3_rresp(axim_ctrl_int[3].rresp),
        .axim_ctrl_3_rvalid(axim_ctrl_int[3].rvalid),
        .axim_ctrl_3_wdata(axim_ctrl_int[3].wdata),
        .axim_ctrl_3_wlast(axim_ctrl_int[3].wlast),
        .axim_ctrl_3_wready(axim_ctrl_int[3].wready),
        .axim_ctrl_3_wstrb(axim_ctrl_int[3].wstrb),
        .axim_ctrl_3_wvalid(axim_ctrl_int[3].wvalid),
        .axis_dyn_in_0_tdata(axis_dyn_in_int[0].tdata),
        .axis_dyn_in_0_tkeep(axis_dyn_in_int[0].tkeep),
        .axis_dyn_in_0_tlast(axis_dyn_in_int[0].tlast),
        .axis_dyn_in_0_tready(axis_dyn_in_int[0].tready),
        .axis_dyn_in_0_tvalid(axis_dyn_in_int[0].tvalid),
        .axis_dyn_out_0_tdata(axis_dyn_out_int[0].tdata),
        .axis_dyn_out_0_tkeep(axis_dyn_out_int[0].tkeep),
        .axis_dyn_out_0_tlast(axis_dyn_out_int[0].tlast),
        .axis_dyn_out_0_tready(axis_dyn_out_int[0].tready),
        .axis_dyn_out_0_tvalid(axis_dyn_out_int[0].tvalid),
        .dsc_bypass_c2h_0_dsc_byp_ctl(xdma_req_int[0].c2h_ctl),
        .dsc_bypass_c2h_0_dsc_byp_dst_addr(xdma_req_int[0].c2h_addr),
        .dsc_bypass_c2h_0_dsc_byp_len(xdma_req_int[0].c2h_len),
        .dsc_bypass_c2h_0_dsc_byp_load(xdma_req_int[0].c2h_valid),
        .dsc_bypass_c2h_0_dsc_byp_ready(xdma_req_int[0].c2h_ready),
        .dsc_bypass_c2h_0_dsc_byp_src_addr(0),
        .dsc_bypass_h2c_0_dsc_byp_ctl(xdma_req_int[0].h2c_ctl),
        .dsc_bypass_h2c_0_dsc_byp_dst_addr(0),
        .dsc_bypass_h2c_0_dsc_byp_len(xdma_req_int[0].h2c_len),
        .dsc_bypass_h2c_0_dsc_byp_load(xdma_req_int[0].h2c_valid),
        .dsc_bypass_h2c_0_dsc_byp_ready(xdma_req_int[0].h2c_ready),
        .dsc_bypass_h2c_0_dsc_byp_src_addr(xdma_req_int[0].h2c_addr),
        .dsc_status_c2h_sts0(xdma_req_int[0].c2h_status),
        .dsc_status_h2c_sts0(xdma_req_int[0].h2c_status),
        .axis_dyn_in_1_tdata(axis_dyn_in_int[1].tdata),
        .axis_dyn_in_1_tkeep(axis_dyn_in_int[1].tkeep),
        .axis_dyn_in_1_tlast(axis_dyn_in_int[1].tlast),
        .axis_dyn_in_1_tready(axis_dyn_in_int[1].tready),
        .axis_dyn_in_1_tvalid(axis_dyn_in_int[1].tvalid),
        .axis_dyn_out_1_tdata(axis_dyn_out_int[1].tdata),
        .axis_dyn_out_1_tkeep(axis_dyn_out_int[1].tkeep),
        .axis_dyn_out_1_tlast(axis_dyn_out_int[1].tlast),
        .axis_dyn_out_1_tready(axis_dyn_out_int[1].tready),
        .axis_dyn_out_1_tvalid(axis_dyn_out_int[1].tvalid),
        .dsc_bypass_c2h_1_dsc_byp_ctl(xdma_req_int[1].c2h_ctl),
        .dsc_bypass_c2h_1_dsc_byp_dst_addr(xdma_req_int[1].c2h_addr),
        .dsc_bypass_c2h_1_dsc_byp_len(xdma_req_int[1].c2h_len),
        .dsc_bypass_c2h_1_dsc_byp_load(xdma_req_int[1].c2h_valid),
        .dsc_bypass_c2h_1_dsc_byp_ready(xdma_req_int[1].c2h_ready),
        .dsc_bypass_c2h_1_dsc_byp_src_addr(0),
        .dsc_bypass_h2c_1_dsc_byp_ctl(xdma_req_int[1].h2c_ctl),
        .dsc_bypass_h2c_1_dsc_byp_dst_addr(0),
        .dsc_bypass_h2c_1_dsc_byp_len(xdma_req_int[1].h2c_len),
        .dsc_bypass_h2c_1_dsc_byp_load(xdma_req_int[1].h2c_valid),
        .dsc_bypass_h2c_1_dsc_byp_ready(xdma_req_int[1].h2c_ready),
        .dsc_bypass_h2c_1_dsc_byp_src_addr(xdma_req_int[1].h2c_addr),
        .dsc_status_c2h_sts1(xdma_req_int[1].c2h_status),
        .dsc_status_h2c_sts1(xdma_req_int[1].h2c_status),
       .pcie_clk_clk_n(pcie_clk_clk_n),
        .pcie_clk_clk_p(pcie_clk_clk_p),
        .pcie_x16_rxn(pcie_x16_rxn),
        .pcie_x16_rxp(pcie_x16_rxp),
        .pcie_x16_txn(pcie_x16_txn),
        .pcie_x16_txp(pcie_x16_txp),
        .perst_n(perst_n),
        .sys_reset(sys_reset),
        .usr_irq(usr_irq),
        .pclk(pclk),
        .presetn(presetn),
        .nclk(nclk),
        .nresetn(nresetn),
        .uclk(uclk),
        .uresetn(uresetn),
        .lckresetn(lckresetn),
        .xclk(xclk),
        .xresetn(xresetn),
        .aclk(aclk),
        .aresetn(aresetn)
    );
	
    // ================-----------------------------------------------------------------
    // STATIC DDR LAYER 
    // ================-----------------------------------------------------------------
    design_ddr inst_int_ddr (
        .c0_ddr4_act_n(c0_ddr4_act_n),
		.c0_ddr4_adr(c0_ddr4_adr),
		.c0_ddr4_ba(c0_ddr4_ba),
		.c0_ddr4_bg(c0_ddr4_bg),
		.c0_ddr4_ck_c(c0_ddr4_ck_c),
		.c0_ddr4_ck_t(c0_ddr4_ck_t),
		.c0_ddr4_cke(c0_ddr4_cke),
		.c0_ddr4_cs_n(c0_ddr4_cs_n),
		.c0_ddr4_dm_n(c0_ddr4_dm_dbi_n),
		.c0_ddr4_dq(c0_ddr4_dq),
		.c0_ddr4_dqs_c(c0_ddr4_dqs_c),
		.c0_ddr4_dqs_t(c0_ddr4_dqs_t),
		.c0_ddr4_odt(c0_ddr4_odt),
		.c0_ddr4_reset_n(c0_ddr4_reset_n),
		.c0_sys_clk_0_clk_n(c0_sys_clk_n),
		.c0_sys_clk_0_clk_p(c0_sys_clk_p),
       .c1_ddr4_act_n(c1_ddr4_act_n),
		.c1_ddr4_adr(c1_ddr4_adr),
		.c1_ddr4_ba(c1_ddr4_ba),
		.c1_ddr4_bg(c1_ddr4_bg),
		.c1_ddr4_ck_c(c1_ddr4_ck_c),
		.c1_ddr4_ck_t(c1_ddr4_ck_t),
		.c1_ddr4_cke(c1_ddr4_cke),
		.c1_ddr4_cs_n(c1_ddr4_cs_n),
		.c1_ddr4_dm_n(c1_ddr4_dm_dbi_n),
		.c1_ddr4_dq(c1_ddr4_dq),
		.c1_ddr4_dqs_c(c1_ddr4_dqs_c),
		.c1_ddr4_dqs_t(c1_ddr4_dqs_t),
		.c1_ddr4_odt(c1_ddr4_odt),
		.c1_ddr4_reset_n(c1_ddr4_reset_n),
		.c1_sys_clk_0_clk_n(c1_sys_clk_n),
		.c1_sys_clk_0_clk_p(c1_sys_clk_p),
        .axi_ddr_in_0_araddr(axi_ddr_in[0].araddr),
        .axi_ddr_in_0_arburst(axi_ddr_in[0].arburst),
        .axi_ddr_in_0_arcache(axi_ddr_in[0].arcache),
        .axi_ddr_in_0_arid(axi_ddr_in[0].arid),
        .axi_ddr_in_0_arlen(axi_ddr_in[0].arlen),
        .axi_ddr_in_0_arlock(axi_ddr_in[0].arlock),
        .axi_ddr_in_0_arprot(axi_ddr_in[0].arprot),
        .axi_ddr_in_0_arqos(axi_ddr_in[0].arqos),
        .axi_ddr_in_0_arready(axi_ddr_in[0].arready),
        .axi_ddr_in_0_arregion(axi_ddr_in[0].arregion),
        .axi_ddr_in_0_arsize(axi_ddr_in[0].arsize),
        .axi_ddr_in_0_arvalid(axi_ddr_in[0].arvalid),
        .axi_ddr_in_0_awaddr(axi_ddr_in[0].awaddr),
        .axi_ddr_in_0_awburst(axi_ddr_in[0].awburst),
        .axi_ddr_in_0_awcache(axi_ddr_in[0].awcache),
        .axi_ddr_in_0_awid(axi_ddr_in[0].awid),
        .axi_ddr_in_0_awlen(axi_ddr_in[0].awlen),
        .axi_ddr_in_0_awlock(axi_ddr_in[0].awlock),
        .axi_ddr_in_0_awprot(axi_ddr_in[0].awprot),
        .axi_ddr_in_0_awqos(axi_ddr_in[0].awqos),
        .axi_ddr_in_0_awready(axi_ddr_in[0].awready),
        .axi_ddr_in_0_awregion(axi_ddr_in[0].awregion),
        .axi_ddr_in_0_awsize(axi_ddr_in[0].awsize),
        .axi_ddr_in_0_awvalid(axi_ddr_in[0].awvalid),
        .axi_ddr_in_0_bid(axi_ddr_in[0].bid),
        .axi_ddr_in_0_bready(axi_ddr_in[0].bready),
        .axi_ddr_in_0_bresp(axi_ddr_in[0].bresp),
        .axi_ddr_in_0_bvalid(axi_ddr_in[0].bvalid),
        .axi_ddr_in_0_rdata(axi_ddr_in[0].rdata),
        .axi_ddr_in_0_rid(axi_ddr_in[0].rid),
        .axi_ddr_in_0_rlast(axi_ddr_in[0].rlast),
        .axi_ddr_in_0_rready(axi_ddr_in[0].rready),
        .axi_ddr_in_0_rresp(axi_ddr_in[0].rresp),
        .axi_ddr_in_0_rvalid(axi_ddr_in[0].rvalid),
        .axi_ddr_in_0_wdata(axi_ddr_in[0].wdata),
        .axi_ddr_in_0_wlast(axi_ddr_in[0].wlast),
        .axi_ddr_in_0_wready(axi_ddr_in[0].wready),
        .axi_ddr_in_0_wstrb(axi_ddr_in[0].wstrb),
        .axi_ddr_in_0_wvalid(axi_ddr_in[0].wvalid),
        .axi_ddr_in_1_araddr(axi_ddr_in[1].araddr),
        .axi_ddr_in_1_arburst(axi_ddr_in[1].arburst),
        .axi_ddr_in_1_arcache(axi_ddr_in[1].arcache),
        .axi_ddr_in_1_arid(axi_ddr_in[1].arid),
        .axi_ddr_in_1_arlen(axi_ddr_in[1].arlen),
        .axi_ddr_in_1_arlock(axi_ddr_in[1].arlock),
        .axi_ddr_in_1_arprot(axi_ddr_in[1].arprot),
        .axi_ddr_in_1_arqos(axi_ddr_in[1].arqos),
        .axi_ddr_in_1_arready(axi_ddr_in[1].arready),
        .axi_ddr_in_1_arregion(axi_ddr_in[1].arregion),
        .axi_ddr_in_1_arsize(axi_ddr_in[1].arsize),
        .axi_ddr_in_1_arvalid(axi_ddr_in[1].arvalid),
        .axi_ddr_in_1_awaddr(axi_ddr_in[1].awaddr),
        .axi_ddr_in_1_awburst(axi_ddr_in[1].awburst),
        .axi_ddr_in_1_awcache(axi_ddr_in[1].awcache),
        .axi_ddr_in_1_awid(axi_ddr_in[1].awid),
        .axi_ddr_in_1_awlen(axi_ddr_in[1].awlen),
        .axi_ddr_in_1_awlock(axi_ddr_in[1].awlock),
        .axi_ddr_in_1_awprot(axi_ddr_in[1].awprot),
        .axi_ddr_in_1_awqos(axi_ddr_in[1].awqos),
        .axi_ddr_in_1_awready(axi_ddr_in[1].awready),
        .axi_ddr_in_1_awregion(axi_ddr_in[1].awregion),
        .axi_ddr_in_1_awsize(axi_ddr_in[1].awsize),
        .axi_ddr_in_1_awvalid(axi_ddr_in[1].awvalid),
        .axi_ddr_in_1_bid(axi_ddr_in[1].bid),
        .axi_ddr_in_1_bready(axi_ddr_in[1].bready),
        .axi_ddr_in_1_bresp(axi_ddr_in[1].bresp),
        .axi_ddr_in_1_bvalid(axi_ddr_in[1].bvalid),
        .axi_ddr_in_1_rdata(axi_ddr_in[1].rdata),
        .axi_ddr_in_1_rid(axi_ddr_in[1].rid),
        .axi_ddr_in_1_rlast(axi_ddr_in[1].rlast),
        .axi_ddr_in_1_rready(axi_ddr_in[1].rready),
        .axi_ddr_in_1_rresp(axi_ddr_in[1].rresp),
        .axi_ddr_in_1_rvalid(axi_ddr_in[1].rvalid),
        .axi_ddr_in_1_wdata(axi_ddr_in[1].wdata),
        .axi_ddr_in_1_wlast(axi_ddr_in[1].wlast),
        .axi_ddr_in_1_wready(axi_ddr_in[1].wready),
        .axi_ddr_in_1_wstrb(axi_ddr_in[1].wstrb),
        .axi_ddr_in_1_wvalid(axi_ddr_in[1].wvalid),
        .axi_ddr_in_2_araddr(axi_ddr_in[2].araddr),
        .axi_ddr_in_2_arburst(axi_ddr_in[2].arburst),
        .axi_ddr_in_2_arcache(axi_ddr_in[2].arcache),
        .axi_ddr_in_2_arid(axi_ddr_in[2].arid),
        .axi_ddr_in_2_arlen(axi_ddr_in[2].arlen),
        .axi_ddr_in_2_arlock(axi_ddr_in[2].arlock),
        .axi_ddr_in_2_arprot(axi_ddr_in[2].arprot),
        .axi_ddr_in_2_arqos(axi_ddr_in[2].arqos),
        .axi_ddr_in_2_arready(axi_ddr_in[2].arready),
        .axi_ddr_in_2_arregion(axi_ddr_in[2].arregion),
        .axi_ddr_in_2_arsize(axi_ddr_in[2].arsize),
        .axi_ddr_in_2_arvalid(axi_ddr_in[2].arvalid),
        .axi_ddr_in_2_awaddr(axi_ddr_in[2].awaddr),
        .axi_ddr_in_2_awburst(axi_ddr_in[2].awburst),
        .axi_ddr_in_2_awcache(axi_ddr_in[2].awcache),
        .axi_ddr_in_2_awid(axi_ddr_in[2].awid),
        .axi_ddr_in_2_awlen(axi_ddr_in[2].awlen),
        .axi_ddr_in_2_awlock(axi_ddr_in[2].awlock),
        .axi_ddr_in_2_awprot(axi_ddr_in[2].awprot),
        .axi_ddr_in_2_awqos(axi_ddr_in[2].awqos),
        .axi_ddr_in_2_awready(axi_ddr_in[2].awready),
        .axi_ddr_in_2_awregion(axi_ddr_in[2].awregion),
        .axi_ddr_in_2_awsize(axi_ddr_in[2].awsize),
        .axi_ddr_in_2_awvalid(axi_ddr_in[2].awvalid),
        .axi_ddr_in_2_bid(axi_ddr_in[2].bid),
        .axi_ddr_in_2_bready(axi_ddr_in[2].bready),
        .axi_ddr_in_2_bresp(axi_ddr_in[2].bresp),
        .axi_ddr_in_2_bvalid(axi_ddr_in[2].bvalid),
        .axi_ddr_in_2_rdata(axi_ddr_in[2].rdata),
        .axi_ddr_in_2_rid(axi_ddr_in[2].rid),
        .axi_ddr_in_2_rlast(axi_ddr_in[2].rlast),
        .axi_ddr_in_2_rready(axi_ddr_in[2].rready),
        .axi_ddr_in_2_rresp(axi_ddr_in[2].rresp),
        .axi_ddr_in_2_rvalid(axi_ddr_in[2].rvalid),
        .axi_ddr_in_2_wdata(axi_ddr_in[2].wdata),
        .axi_ddr_in_2_wlast(axi_ddr_in[2].wlast),
        .axi_ddr_in_2_wready(axi_ddr_in[2].wready),
        .axi_ddr_in_2_wstrb(axi_ddr_in[2].wstrb),
        .axi_ddr_in_2_wvalid(axi_ddr_in[2].wvalid),
        .axi_ddr_in_3_araddr(axi_ddr_in[3].araddr),
        .axi_ddr_in_3_arburst(axi_ddr_in[3].arburst),
        .axi_ddr_in_3_arcache(axi_ddr_in[3].arcache),
        .axi_ddr_in_3_arid(axi_ddr_in[3].arid),
        .axi_ddr_in_3_arlen(axi_ddr_in[3].arlen),
        .axi_ddr_in_3_arlock(axi_ddr_in[3].arlock),
        .axi_ddr_in_3_arprot(axi_ddr_in[3].arprot),
        .axi_ddr_in_3_arqos(axi_ddr_in[3].arqos),
        .axi_ddr_in_3_arready(axi_ddr_in[3].arready),
        .axi_ddr_in_3_arregion(axi_ddr_in[3].arregion),
        .axi_ddr_in_3_arsize(axi_ddr_in[3].arsize),
        .axi_ddr_in_3_arvalid(axi_ddr_in[3].arvalid),
        .axi_ddr_in_3_awaddr(axi_ddr_in[3].awaddr),
        .axi_ddr_in_3_awburst(axi_ddr_in[3].awburst),
        .axi_ddr_in_3_awcache(axi_ddr_in[3].awcache),
        .axi_ddr_in_3_awid(axi_ddr_in[3].awid),
        .axi_ddr_in_3_awlen(axi_ddr_in[3].awlen),
        .axi_ddr_in_3_awlock(axi_ddr_in[3].awlock),
        .axi_ddr_in_3_awprot(axi_ddr_in[3].awprot),
        .axi_ddr_in_3_awqos(axi_ddr_in[3].awqos),
        .axi_ddr_in_3_awready(axi_ddr_in[3].awready),
        .axi_ddr_in_3_awregion(axi_ddr_in[3].awregion),
        .axi_ddr_in_3_awsize(axi_ddr_in[3].awsize),
        .axi_ddr_in_3_awvalid(axi_ddr_in[3].awvalid),
        .axi_ddr_in_3_bid(axi_ddr_in[3].bid),
        .axi_ddr_in_3_bready(axi_ddr_in[3].bready),
        .axi_ddr_in_3_bresp(axi_ddr_in[3].bresp),
        .axi_ddr_in_3_bvalid(axi_ddr_in[3].bvalid),
        .axi_ddr_in_3_rdata(axi_ddr_in[3].rdata),
        .axi_ddr_in_3_rid(axi_ddr_in[3].rid),
        .axi_ddr_in_3_rlast(axi_ddr_in[3].rlast),
        .axi_ddr_in_3_rready(axi_ddr_in[3].rready),
        .axi_ddr_in_3_rresp(axi_ddr_in[3].rresp),
        .axi_ddr_in_3_rvalid(axi_ddr_in[3].rvalid),
        .axi_ddr_in_3_wdata(axi_ddr_in[3].wdata),
        .axi_ddr_in_3_wlast(axi_ddr_in[3].wlast),
        .axi_ddr_in_3_wready(axi_ddr_in[3].wready),
        .axi_ddr_in_3_wstrb(axi_ddr_in[3].wstrb),
        .axi_ddr_in_3_wvalid(axi_ddr_in[3].wvalid),
        .axi_ddr_in_4_araddr(axi_ddr_in[4].araddr),
        .axi_ddr_in_4_arburst(axi_ddr_in[4].arburst),
        .axi_ddr_in_4_arcache(axi_ddr_in[4].arcache),
        .axi_ddr_in_4_arid(axi_ddr_in[4].arid),
        .axi_ddr_in_4_arlen(axi_ddr_in[4].arlen),
        .axi_ddr_in_4_arlock(axi_ddr_in[4].arlock),
        .axi_ddr_in_4_arprot(axi_ddr_in[4].arprot),
        .axi_ddr_in_4_arqos(axi_ddr_in[4].arqos),
        .axi_ddr_in_4_arready(axi_ddr_in[4].arready),
        .axi_ddr_in_4_arregion(axi_ddr_in[4].arregion),
        .axi_ddr_in_4_arsize(axi_ddr_in[4].arsize),
        .axi_ddr_in_4_arvalid(axi_ddr_in[4].arvalid),
        .axi_ddr_in_4_awaddr(axi_ddr_in[4].awaddr),
        .axi_ddr_in_4_awburst(axi_ddr_in[4].awburst),
        .axi_ddr_in_4_awcache(axi_ddr_in[4].awcache),
        .axi_ddr_in_4_awid(axi_ddr_in[4].awid),
        .axi_ddr_in_4_awlen(axi_ddr_in[4].awlen),
        .axi_ddr_in_4_awlock(axi_ddr_in[4].awlock),
        .axi_ddr_in_4_awprot(axi_ddr_in[4].awprot),
        .axi_ddr_in_4_awqos(axi_ddr_in[4].awqos),
        .axi_ddr_in_4_awready(axi_ddr_in[4].awready),
        .axi_ddr_in_4_awregion(axi_ddr_in[4].awregion),
        .axi_ddr_in_4_awsize(axi_ddr_in[4].awsize),
        .axi_ddr_in_4_awvalid(axi_ddr_in[4].awvalid),
        .axi_ddr_in_4_bid(axi_ddr_in[4].bid),
        .axi_ddr_in_4_bready(axi_ddr_in[4].bready),
        .axi_ddr_in_4_bresp(axi_ddr_in[4].bresp),
        .axi_ddr_in_4_bvalid(axi_ddr_in[4].bvalid),
        .axi_ddr_in_4_rdata(axi_ddr_in[4].rdata),
        .axi_ddr_in_4_rid(axi_ddr_in[4].rid),
        .axi_ddr_in_4_rlast(axi_ddr_in[4].rlast),
        .axi_ddr_in_4_rready(axi_ddr_in[4].rready),
        .axi_ddr_in_4_rresp(axi_ddr_in[4].rresp),
        .axi_ddr_in_4_rvalid(axi_ddr_in[4].rvalid),
        .axi_ddr_in_4_wdata(axi_ddr_in[4].wdata),
        .axi_ddr_in_4_wlast(axi_ddr_in[4].wlast),
        .axi_ddr_in_4_wready(axi_ddr_in[4].wready),
        .axi_ddr_in_4_wstrb(axi_ddr_in[4].wstrb),
        .axi_ddr_in_4_wvalid(axi_ddr_in[4].wvalid),
        .sys_reset(sys_reset),
        .aclk(aclk),
        .aresetn(aresetn)
	);
	

    // ================-----------------------------------------------------------------
    // I/O AND BOARD SPECIFIC
    // ================-----------------------------------------------------------------
    IBUF rst_IBUF_inst (
		.O(sys_reset), // Buffer output
		.I(sys_reset_nb) // Buffer input (connect directly to top-level port)
	);

	IBUF perst_n_IBUF_inst (
			.O(perst_n),
			.I(perst_n_nb)
	);
    // XDMA 
    for(genvar i = 0; i < N_CHAN; i++) begin
        xdma_assign inst_xdma_assign (
            .s_dma_rd(dma_rd_req_int[i]), 
            .s_dma_wr(dma_wr_req_int[i]), 
            .m_xdma(xdma_req_int[i])
        );
    end

    // ================-----------------------------------------------------------------
    // SHELL
    // ================-----------------------------------------------------------------
    `include "top_shell.svh"

endmodule